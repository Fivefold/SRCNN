library ieee;
use ieee.std_logic_1164.all;

package config_pkg is
    constant IMG_WIDTH_MAX : natural := 300;
    constant IMG_HEIGHT_MAX : natural := 300;
    constant KERNELSIZE_MAX : natural := 9;
end package;